

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
J7NzBcIPSWRzNRBarceM2DFHC3vA1ZU4yTRCkS41yz/xrpSO7Qc33e0okpNQhgZ1WwudCAhttNPu
UUOY4OF8tA==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Zjtm307Ykxkd4bcBuTA01oTvGN3JCkUPJhrFaZvF1u1HdlVFL+CdgH/mJMTpuKq/qLIcq9qu3K56
aAo4vtj7plpHhfzYfrC5hEYegM9+/OpjKHnBFRzqoeYyn42c2JS7evIoyfrpPgu7EcCdJyFSiE90
L3ZI/Mx69e3ZbOxIolg=


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2014_03", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
c6x6FARdruHUtc5Z1Bu8NyKc9zznCeoLEIOsYA3WKEt+78TuKZhnqjbErSudJR5nXQkK5iZT3bJX
h5isz6jHdM8l1U2AZnpeP3XOM3yexU3j2NNeR9v82jU/6+Y8zN/d/Xdx5H3uFhfc1eAgw/JLoXZy
qe9j/EbUq0+T16ZC/5FzefQSWpQbjCSTeBGCqwiKuLrdo5c8mO4xqxdC/bp5cokzEzmL7hAHMS86
tscXjBfVNX6QvywuuiRqVOuRbxRJD+jbVDrhw3m0T+1XEDD8Osn4FgHAhPcMgihajKOIwLKeeg8I
Gcy10KwpwspgrD5ZvYNSnvo50ZV8vGkCT8soFA==


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
3h2iw8H8fgU0xT2ADEB3q3xK0+YRgmH54AXa+fK7z+LUk7phjT46ArfJriTIn2n5qKQvEY1IIHPC
X/nrcuIpLrY2Cd06ll/zx5oTBRNA7qmTitbIbAFocsxp3rqgEQJ+nL1VQlbHwKRT0o5rS7c0+L4o
1vz96XsuzmXTgFA5mFU=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC08_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
fIpPQTsksNLtapsSf2P9IQqpskDBe39wHYkbzAcYN+nyuus133ITXmDqXJd5a5nRnXn0gjSEMvBx
2D/GrX4TGxAGWVRnNqheKqM1EXeIhv93SPKdhlwrMblHE/Wfr7QhjkLKS5JQoTXFhGNqub7KiP44
ZmIIxkF19gJkPYtHlhItavED6C25/KjN6mBIDCmo5gqf1To24xOOGiOAtJ1xjrChUhd0zzz7oeHE
7nZbX36KvSBoWIMY/+KJGjnib/IeX8NClT8a5gcqg0CoqVJ3sR/jUkzuVBU+e9cfHk9VB0h5yYYB
3qi4omCKRf1zpWbhiCizjpB7O9Kjg02J9iigQw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 13456)
`protect data_block
YaQlFgHnmPqBND6VPuNTBO57qZxufz5s+oBbyWe6XfkROEu+OvlfOSRyGwz3342t4zfM9Idc7cfY
cs9oEJFztksFWgPghhtaUhCt5neSOCMEsp/Q7vKDZbNcE+If0QXYm9309yENaqDRfIcbWQir2WSf
WCgeXSt+HPCDkJ87qd94z4E4erNWUWekb8bxCL3LKZI7HCHOyhJUedXkGf6JLBRmsBZ9GbnC7XLX
d0u5qCK/xeDJcMsgZ4nLH78H7ibHq4hxdJFkdfoC5BbgiE4PUddiY6SZIn/oIKsAriTRGCCCmra9
6env1sARe8CiGv5el7aW2m+R//EgMsIEFCkjUBbnqxknSwenWh2T8RLyS0e9lqOgGm0pDKCxjAaW
OtpQgXcoLLfB3zaJNaCJRH9Od+NooyFs6rX3pkhZ36zXiuSndmLL3MJhxJHfR3wFWcg4tzqNT2a2
3DMGHcHvLC0B0bSoM1LH/Y/rGyy6frPCzO5fVlzRou1aCt9ivn+gasAT3A+9TPoFzAEZwDaxxBIC
iNK+G3fh+4trJcBLIYA5PV/oQpdHyLQWM7soLZMpNbCRZweMPLMANG47VC5JsK8NsqlJEhmP5CmN
Y00UF2qwTASLbsVI15JM9fKoxhgEzS6OfUrn+/WqWwb8c8E16XAKViKFgkf4ZZp60cVWfgj1D5Wc
lO8zvROdBrgzDq61Z8RxY6YVSKeBswJqYuavt/eO0ksCrA8NuQaKBEc1Dv2v6p2WRpt9TDlrHLOe
xTNerFbAC6k2ZPjoOiFnmEnv/j3mp1ldHgXP4dVbiKWgC+Y8s2LtY+mYOk/LAVhMSiIvsG8wzYK/
Rw1r16ft1dmht2hIDTn/75fJRsu+BRxXqe3EljYnX8sOMWWgVk11xW2aVELJsdGjlyPdV4ZXDN2m
Q8qm7vIxNTZkN8PvtdF0eUFMBmhwlkOwcp5nUFWMTCcOgHCi/vTQ8F1QpxqrpI6T1TGRmvxlWe2Q
aKW96Q3fRMb4cVnLhgdz1+rzFbVIpFjFSlwjIMFhuPCvNP8JzVvi2GdNCncHw0JnNNhEFqYXBcbo
tkph1BLIRQP6Lu4zpkxymVk0xlUF76/QNrmI9zWDTdKzzC1P0nB93b3MSDR3SE9A7634Mod7/CxX
19KbtXMwBotwHjP3fZIuuTpeTEYQOZ+cMP0fJa+NqoN0yCm3DcRO62WxOBKNGTrz0ae6VA4Q9xxe
8JRtceq+T2B5NQIg1Al72WzpXwkKU1lOSRt4cjAu/NwxJoKvXo7VDt9WzdbPBtKqkWDuDWoRvD/o
nByrePDyJll0SyuLacciQDB3X6YIQPtzgSsTEGB063RgqsbVsZVaahH3kM5WUemu/GWtgPg1YI7V
1IVwXfUZYkBQ16IefCOHX9vEYjHoeWpMhya7vcZ1Vt++BWz+1W33xMKgktBPVn91L+ei9sG5Jwww
CJp0lqiaqmK7we9o+tf9xtI6UpeyDDRXptS48p01EHI6W5vP+7G9DaxtKWYL+JsAQkZAOVOlTSW9
NHPcwrFXjiRCHnJVIFTgo1n/Wh0vVeO9Okvq0D6KXhXTUrOqhC7SYx0rt3dsyVlVsfKAiHX2hG3n
erXwBrB70N0HMMTNucKo9h1YlT19dmzxun71KpGlhc5jiipW1hbGAw82GE3Zfka9ovPd9IuXDqIq
5twpg63CTl9WAQIcs8yJFuCzWBs98jqRDX1J2CCIFMPHbY+LAw0VGGnaARfk55XjAMoW9YdX4kyw
6Hus7nw96gVJ6v6jazAgac9gbwWt5ebNGI9LAa+YOwnbh9+zJ11xwZsADOizqmZoqQuJfObD3rzx
GX7qQKyj8u6rqy/+s+ktXhKiPepO+KT1/vlO4t03w2D7PaOgfsoPiL4V44pB56lisWQnCpfHg7a6
V1fpe6vqMD8U74pL8BRLeePEaxyIN0qbYTw90EXMWeOmqz7gBRBnOHiz4tmJs6YBxH/FSSZETZ08
OYy99A/mKHEbxmNaa4z3IzGNfa+G8tX2/pKDKEJnGD53QKKElEUQmHSQj20FC+G0DQFlok2Aq46D
5C40v/+y2CKK0IIbOV7ZuuwxvLjeYGpND97YrhFRa5FVcvMNj5cL9Fxv7A1UCrmFB/49XDWG2lZ7
PSk9Non83DWlDJtdeFqM4SlWnwEZ15oPnCgE11MF8g8CaBx5jzCS1l+sMjgImYJNRI8SBBQfAp1v
7pfETKn8fAt5RJkJcG9G2FrAz+d79COm5SNEGEyuriw3SkG3iA3L/2OksLzkM6aF+UhPPn/8cDFf
/siiuQ1FEY1JobuwcxMtSgLMCI40VNkTeM36lu83WbJgpWgn3wN33x1TM0kbFmEltasavAigFUQF
B9xRZd4oUeg1lthJ/qtqkUA2y2Hlppmy2Fm1xzn7NC31c2c41YHQsRJWxVoJcnUqFHzRFcbc2u6u
Bs3WeYYY1VKzm8Plre+Azi0/q+W6BnU4WeTyNfSsUrGHgWe/Pmxo8H3aXB8biwUY7CtapLQXbynZ
7c+Fgr5AfF80H5pyBB/b9Nj/h05JgapLy54SNQzbfbZEJQrD5pjHqoYC9sEHokUcwV3yxNt8Uk1A
AZsQTdMjiDVNHx/dUv4hwJVOO+MjrWPx1gk6FFJddA7mfFfPqCfm4VzeAGGRN95NKUBoARVeO1Gs
xAhXaGEYg7Ee9z2xrtAu56efD5bYuudVW94FC75nYNp5xdFz3NMNiwygt06uwZI/aXp0eky7fM97
KkyzsSvY3wePhlQ2xlwdkSknkXBN1X+oS8Y1lr84Pz2EJ1lhg0P11X1rVqJfPV0s7qiYVcl23oBJ
hWHrnqvs3Z2d0xNvkav7vnHbP0pcml8hVl67z6tzEsbPgaDpNvZUwt/YWqRB38GmngJF49kr3ZvO
ayRK7otIQs60Xh/PO/Ja6wj1F6g5+SGMP0S5J0u2uz2pD+1LAga1rMnhTGN9/OkB/08/UZAuQvyx
6sBd9SC3s3r1DaV3jmP+8zhCmLv3c7zanKBu+y5BnwXeUCbtKhU95bPB5h+cX/+Fen1ze0llrYFd
+ubLoDlbIOBuY50sCBMfwX5neU4XllWGjRDAgacG8WFSmsNwKy75mRGD3dDmMVDQ1+en8PjBI0Kp
5KrpJPjm6MB9kLNp+nYQd3OeM+M9t9yGF+kwwfhInXgBr7m32zei/JDbKVG9UvkwIprO215OYoWO
UP4fPCnWRlHZ3dA7tyBeYzt0D90STPK0p+htYtRydrrpWXR4rvRal8rau+mpc8mjiccIwZWKemjS
85+2p3OXeZjxbUKgiUGPSxC+tNPdBwXKZ6dnOwBsAYPACHkqtOUpFxdDjqO1yJnFowZVODTYYBq0
va3WiEBEalKIsiMS5hA6x3f/hwW1mO+xSG/+ir7MlAh8VheUVVErDtxs4Us3esanqHUOHLhxgndG
VSWlmfSIk5MQwhLp2Ye9n6HviSdZFc8CM1JC2to0aF3GXjlbqH6ZzvwTwtSK5/XKX4ZbArr4nz+c
cDDpX41hNXwrnX7eaFeFo5AI5kj0EfGFuMZZWuPH6s6i5CWwBXesKP4+q6n/QrnX+vYTYZFuDXYx
eEenXk1ZadnT7HJFM57k7/lOXFPMntCkCHDBFCIEW2P6WYzRgqND2P7K2uJCbgjFBpEe+VnaPyqN
Tz2fcEAlP6OGomGBC5y6Erc6l2CoxWYEos5+1AXXKjbOO8Hc2HbrtfSLR+m2Jh92c7UQ4MRVa0/9
L7Tlm0p+Si5rzE6b7qF1Bhwyh8j/tDRodrcNdFCn9dlc5tO26xCBLVO7kVO6OVjDojK1U1Ew1/N/
/1LnnzprjhZSlm+ipkKWqXFmOoWxCGodeF9Jj2DHnXHrhxkq0TMIvxPXUFNxwI4Hi2PZ2QH2D6hn
166mmQK2Y5SqR9NIJIfrL92V1xQtpr44GGGdIC1TOwl4xUKOy6n3tMLl4fa2FOXjKhTZwmwUmY9l
LaiMZm0FF0Lt1Nqv2PVy0eKj/wImdyeTm+07lTbM4kT2nz3+Xa6E1fCpltfyeNpO9CApYJe8UifE
PL/fYa/3wS0XHRcxWRVwzlP0UE13w84OevNpZ1J5hvQWJTeL3GClwjPIYXihtvOJtFFMrEkCDqU4
UF3uUYgnTe32Xkp0pi7+0tunR5xiWRLZmFY0oLf4ci2OGOKef7l+zUexMOiAwMeDfRM+ul2z/j4K
fbVPWAx8rW5wxrJYP9voclnKF4HMkGGgSYyjjQ0nIabQzYUrwU9Z7zVh0WCpJr4s153trymqEmCn
xJ5krSpYqDgpTnSDHJmpOa/cDuA0/QqDhgWfTa36uF9dM17gUAgZsjT3rF44x9yFCTd0Ko5/e56E
ydj167nxsSlVCx93j9t5TTjN40dTXP0ayVIHyGb99SbKzrbBRDQa/rxcOnQA5jD8XnrzELq9R5IK
cJeumCoh41ErQoedOU4rIsGiTSnYK6bur/rDd52hztyqDZaj13ZafSURDcQhXQEeUxhSzSqFS0DD
5dSVIGvgb3UgZajxzTIe8pF7o1hzf4LY0ZwZyYVOfmmDaEy6liByADKjsY7LgnBy3AkCuyu6bBau
svvF2BOiMEOGUQqDkpm8CCv+C1lQSScvGZ6acjYFlPYokHTQnVPr6hppXeUy+HJL199wapC7sWcn
g9mO8Ujt4XX+F+vCzYNllU/P5w7B4FXm1RXjhzJznWN+jY9adbezJ8xybgrX9Rb1sqvIu+4xLr3f
dS1GPz0xjlbhgEGhubYGNl7zUZxPG5qHRUca2qQbkRp2Vw9hi1FYWd0plW33OBntS4rv5kiszEq+
JTQI6dJgsGlwW8CxesmuwtOK2cm2MTVleJQvNH2U2O8FZhiC4CaJAIdcev6hMGwEgw4tTYwTXgb4
IwUE1r8HSmwm0vYhq5KV2NyrvH3OkD6DZ2apOZlqSRnGcYfX3k99er9Ahhkn0OjdVktd3x4j8eiR
YX2937yQ2sQ4Eyci61+zyH3cbAkK4XZFlErsNPpjUKtKYRJJKTx/7eZt8cewdP02lp1l9gdV+ajS
qcKc6RDJugBSveMS+RrYuq2d2RU0MZQKYvyZ4dA6lCyJ9GXgqtTyHz8Gd9DPhbAibLLsqlZNg9tg
5KJlN45lFy9d1aJuTRu09qYQEo/g7Wg7iKLIob/CImBcTbM3iqkZZlN6sDhdHnSB1gawQy9vCloK
ASCeyiPTwv6/XFasT/coEcOAcAC46IGZ3VJ9AbhS/mI/mhRBdlVkYcWB+ngB3SLmZKepUFw6FJoe
k8GG5KtFmDPvPlpWMJ6Wtp7CIXQD5OOcTPK/l2nv3KVXqiOGzx4s6QPMqdks5rYnDYAhNoa/i7iP
u3ZkoWMiU94SH9uzvusFXTF8xzDXPtQ0l6nJPsA2w8xQoalAy9G9ESxUw8UBpZGi9Cx6aKueBvjG
gy8U8lOqvECpxW7k5563kOUV90qEZH/RFJVHBMZzl17/6ScxoRULCAdDQmT/T9ShdnPaqSGeQrOB
QXbbnsw9bmmPsl0W0oNHIUhZtlvdxydMdL+tzxGL03my9Ln+MhCz0FUh8XXMWUMPuCbrM1Hn4Zv6
VUlRY2UeFAg6w92ENH2ZeS+cQjFoGExRV5Wd9KcHRJtFFXCy2eLxJLrQ1KQLsXGt25pv8c2Z0qxD
JVrDjB8MmCgmVl/IcyNQLB+RPpSU573NXrJWCgKbDx1+cbA0LXZLcXdRlHtKzJrU4DKYLjW4cg9Y
+u4t5pb3M9bBWXYRjen0WmWD6PfZeK759aQrGUiEXZvsZaJCIOeCxPlEaiCuoTC0aJxkvktpIvw8
7nP8ecckjvZeH9CHC4e2fVADl1R7rJQuZcHAzbTOUrixy2IlpQVWdxh9yJ+OtRoSxQSISQYbSiY1
6j0oH7kNpMJkd7LNGulAZ6U21xTMFnflu/FdiwAdkMYKRUPwglP1nJP2D3Vplxh4fF0whbj1yGRj
bVKv6SW0DPU/S1P/qlkX7NACRsApEskBwbETsiVsQt+jQfrp/dKuA8flYSSWosffTAA17MVa1zxB
ZP8PWLGozlfnU+QVTONwC0/RPz6D4xfiYcjeOTQbNOlzYyKjFq5p905/8/w3CH4N/u667QymA581
8Xqf2fhPF1syT0oSJp5U2dj11lV0TlQQ1CtKEg5xoQ+9R3iV4f7xjJKgEajVRDnDSTVD1iB4WwiQ
cNCGzKvrw1lEpl1IlIU9xqYP3wOPHEcqz6bL33UnNCG9OCNJWcQ44J3Jb6pGULjpnwD3S/ZZRK/o
v9XWAjQ8ir7WafM9gpA9JY6mOvLKCCBfJm4iuzUwZ54u3C3RMJ1kZRd2wXzecT3r7gfzWZrOtg9c
2/P/QKqVrgrp4JwJmZY33n6qLK5/K/CTtC97NrRw7BeippVTFvpuQcm7wsHmP4XgAwst0iqIHltO
caRTLHhsxJ1dhApZxz+L289+CjnK3aHosU+2mxz/I3FPUGQuGts7tclYGbeTlSub/wdYrW7XMBoJ
QoYBPRVcmOacNCitbS8hVDiftyX+/A26iIlk4NqXoVeC89PY/QBTX6Ufqmp4gii0gQxtMqYm3A71
CNWL/rLiIgg/YsVoJ7l/e4WxY1qvFpp/H1vciDOFeAdfRKo5b8zcOfH9DGoBB5xZSfQjKVab59uI
Mfq9xQbdN3xkTUEFdlfsyFnJcGdHk6b37Sqx8F0P8NOlByyUFmU7Br0PK544ZfdHAo/4NntUnQ8Z
lZZCK7J1rIp5KVy0tdGf3IVrxRydQSCIpT2THRVeKhXNUcAHPJ6KeSJDGvJLbzZsuJm0TGIxHH2o
ZvJ/orAYK3MDQOQ0LigGtXMGLJ+gEi2LTSZOMuu7O2TTpYNr9FmdvTGw6uJpGkaHAABtRfeJCirA
5TXdWv1NZKfyiGqdAoxw0lmcDOJE5Jr9v9lqDNVvtSKgch/K0mrPSTg8IcfLBs3SnFf07z/beLe1
Cxuqo+Ggz62hwMz9yp3UO874lUjPdPN5c2xL2NEpacF6VejS1fLlsLjUhYjgU9UGUFkNnZLFcAuJ
xfmgY3tw+jbkRbAAFBMTsw0+mzJYDYYT8cW3K5hTIG70KIiajmjR7N7eQofudaM8CpAWSw45D7yY
0ZTYGYOsspuGH9W+WOfCyGCbnr2UpzpH0Gg3UykXQle6cRF8DyRKfaS01F0QwI0RgE0M9Th/3EYp
AWpdB8mKaoP14L1M4+ezUyj03mDBvaaQuSmYcJIAJFOL1ccbqIme0kdks5O2wP4kTEMflYht4NGf
rgwbzDSj67ZT52JBcKfnBaqf9vDBlVMOoPUvLkDcSBVepb0LqNj8sJsYoDox613FrBoPyDKiWvsf
lgNhtaOQgdckgZk07UAPcarLYu23twthEIU50q8qY0Gb+RCbIkPjkG5hyaxrOw0mJfbRmIDIbsod
Q7tSEqcxtH0Ba7kXPWcPsWpECcWBDmzflP1/rRI5YUEQMwuhMwC9FCR5Gke/HkGXz+zZ25acRl0C
jnXfiayh6kvE2Kcb1rVu4FnoHrtT4ABOZULI97+Wy60LrvFLeZTWeQ9wvPuRYkfYTKlMSdSxofU/
CWhXDoUbUgH/BK/icUl2dlvrJWHHcChpK5CIHFT30lXTXlnx0babf/OyUI3p3pARCtPktcBdqS3X
zkhzDYp3vy4JFXdwebdVHb1txfirUM+QBIawMhhNz3/zny5TAuE7uHD+wjJGzfePzFLzH9qgmMVi
nOoJy88qBLkNJNWHHUqumwkH7DHMWsLeIsd5VVbe5rfC5G8ttiS4TlRPoNXsDMN2dxejYhgTfJVY
gzHw6kRfnYx1FxK4g6fdjO7wdL/J/HVfRzVOh6SqhctObn9qZPSn3hXivYy+BsHctKh+4ClMpAEF
JSyixhGygvBtf5Lgg934VpjalQ1YgUbmHQct1AnRsy4bcusiVHfFpK/yHxDHZGQVozwEsjkbSOyk
aS1WGD+eTEQ0obSlFDbFYhigzWqeWQhxAgrXYPmpKEP4iii8qp3AfNA7RZE+Tow5rhlug72ADtF1
58H/l+f8gIPWOtejmlzKzdw14DL7Gl9E3fEY22C9CwCcgq+FzYD/mXJ5ZZP9ZIWPTOdddsoR2FVJ
z7qXFmg4u+/lYTV91TmbqMpopEJ/mMsDRT4ZTU5zkL1+8o5yPE1swsSUEu2pHpjYNUw9vXHjRU1Z
NRMmAHaQCWXQiZy6dk3rriEiwA5SSFIQBNtaWTlKpD6mVSIbri5/8jbimB/ecMSnp7AJi5LwnO1R
jpka6tyR0RU12iHIbJipSeuh46NAwqYlLLr6m5456cbIpITHs4jyonN60T1cbWIjPfO0asak6l/v
Nptc/m3lHlvDd2sjYb9AorV5hdGyYAFlyUpr0HbSs8ABdTN+a7Ec2KqUVQC/azqON3f+tyRRJUY1
7l8D5pHXdjVwGNiiDFisNfQz2NHYJwrFIPXJEWZmNk6t92kSX24OaLdjoY9qIRt5jnXSP9gZ5Tkt
NQox7c6akdRYG/tJRCRJM9FINicHdwqqKi658sQvdQB5YobNw5gytNSgjwSZCJMp42EHam+r/lKc
Ud6YtE7RQPaoF7KkrFhmBVoCC81Cad43zHZrW559VYAQrZkvVEWNY548UB8cCKuEQ60/8EAZX8Fu
Ko4dzwXmU0vNa1VOldMo/aS9OecqB8DfQL4HKDhiP5kMz/WH8RnoAPVlPRfwa9Ok2efYw1ORzG0e
raXO+EWcwwMbJxFBIxIhW/YzsDFtKXNWyFKqduy+zVX728YWAzBkY/yGEXU8W8vK1N0r+1E9mn2y
gLHYVOXGJMIv6ko0OC+3Vku4ldAp5LPWwUyEsKsd/Ab+sUO0wkOil4M5WPXNhNZ5nurHj/IjPZgL
5p1xO2Xpu9Baj436SFSbuG8qB6+FcPk2CBDi81+Oo+DzgPbK2pIDrDoaLZ/p4qdjBZMn/JE/r3Ez
59PxH8MW+2NYbPy0ndDWGAsP3HwSYIztE0CYkozz7oXtQp4uipXkci01yti6s5Paw92Br7eenhWn
DfgjyYM5pBdA0g3nyuetJz0kJwOxe45z6sHFi3/NjXkr4Xd5TqQp+LhseR3MCSkoeAStm5O3bsxo
adQlxSxzB21B1E0i3SKCmoJ64osdgru8zunOjaELR0T1NEMk2HsM9+MYUENme1wpl/dkQra2LFuO
9ok3E8Fxm/xkQELo73NYB8MxmccBG+OtMlDQonN9b8cWMVk6bMNmgF/vU37BuFhgpbhvWbqnHSCI
/nsBq/yOp4tqiFhcOg7/yRPBa0E7MaSdebzXKtgFDSikIp9a5/xw0g77BzCRKcsxBgPfRzO20x3p
74GOtO5wsKLlmfoQfk5SzsuT1bVzVW8eUFJQAq1I51x2QLRO+bOlbmb/APgylZXBVvLcUc2mFLJP
82pCIsfrtTCz/jJWSaDHFkYBoiuFWBp9vNY/4Sfw2tgz2USBx9psR/rk+X9j9jQXcwQxWwfV6oVb
+iHyllsWfcN2dqL68VJjfWUg1v0Bsh16LlRUer4CWbL4c+sCgJq7tsmX4izk59e0Xhr7hOmE0U8J
03QEa/5+HmQh69f+Wb/eD7hDXKYOtF3dXWvvFfhwh0HotRda4qYvlAjskNoFmbJW8rM51MYyjmYg
iDvI1ybQLxBisVcmjVcM1lQZKVwCH/UetgNhJ6IIKoR2hmpbYHdcKk6gaI230p1gr7VSOQrLy7h0
7FY+Vb+tkFStTDjqaVYAQQw5vc//rmZCcH72UYpfK/HylGMSA+qX+tAbivv34iiN7PC4XT0Y7Nzv
bSHH+3EENnMB2+uRcckW6Y46QPejX1tlIlunHAb0tgUjjL03SR88Beb4LIcMwObi63TljvgIVkwX
ecAXjlALJFOozhNg36qkkDNUoEleuOMrpVkekEeH1LlitcOeH68THd2x+y+y0CBK0a3uqe28dFYh
R5iaEdPJKTBcwIyN7Fqr6nKKHdaAbZEnEa5D25WNWOLRMOlQ7SPNTRSy8EOf10d7pQck13Mhj0du
gOpdDB8IjBAZ+3MXeRMEp9G2R4mg3MC3x+1EgtTSpgqlo66N4iotGGZdua1o0t0+nprlm8DV7MBq
hmNvxMEYq4zq3WN84YImj6O3RjnqD9OpqQjHksH0OVX0aeIVsa3is0gPN/qKaLSyJy8x5TRAYj0Y
ULgYHfr9HinlvPdjGrv+KlO+LFQo6PMKLdjJdxYL+wOhHE77btKwffwg6FrRoXLmAgX7b3nAMqt8
GZTO+8fgqdT16YWJ+Toq5Uv3VvwuQQY6y/xLPGuRi9Suzr2XpMcKn0jpEY37HLkKS2j+RezLvwGo
OL96cD55wRejOF93qAXhlzOAU7d3bIjdCdFI/gjvsPpSZkSCj76ZMz5odJr3mtjeDPgpgHVL0aXI
523fYSl37No18TVomZJNlPxi9uaVWnlghEWi+fkBxiCXITKqQ6OUdC1GR2ca/FroYEuoWhWIXaVK
4VVssd4yOcrl8ZLxi/0dD3/UqOajTqnRbIcXtjN6Y3M6SglBBCbMwcK08KTdsrdWzJbe5d4XNA1l
9SMjtbrjICheBmOaDdx1meOLHbkAO+CrVXfHGL/g5AWqL7ckrPPQKEmdtXMvyLeKzO2ChV5nCNGS
lavfgvrxvkngGRoPXyD2NuJJwDfzmTdGm4ssQ04tz+CQ5TV2dJXOzUDoRX8cyTe63z62VSxJlcO2
hcElz0wC7ThY9asIg/LKJqKsOn5iAPzvp8xoEWVaP4ud9+I1NkH0Sl4h7Fe/LeIg2y4ZiQJSOmHd
X/X1IzkDMTv1zplxPOgQ826WJsgf8bFCPALvp3nt5qECjMI4RDMw70EUKZXRKY6dFnMDqgRjzVbF
nEmb8N4SJ0sMAilrln5KxQum4yLM8w2LWUfbtr1pUCRfRSewN8lpd8mZsAKVKYa52p91aGIKOZbu
+xZ/OZaZt0nTFex5OlwiJnD4QWiBUf5VMjTu1RD2SpYb3pCqV+onAYSIEBjYp7VAsjqiMuc9mIzP
o6gkJipCfQ75jAku/US2x7CXiMIffFS6ne7MAt/WrqEoROgI8LtPha4rB7ySWDg6wODmWUNQDzwf
R1rJAmqOnsOoSXXTKn9dHdinupF+tVEOkr9J15wN8uERqdUU/xQ3LW1Tas1pS+N3rbZ8U9/Y+/d1
6i5Z3Q754SxKsnb8wjsB8mFqZhgsYckVg7G0Cv3VrKX2+nEMHwe7k0XYDHD0lwMW4wTHax/O7zc+
CP0UhYsS4YzCZB0v/aiKfrAdWwWrDL6yijnA0vt4s5cIhaszXTA7tDzS1SOa/Qpm1X86kJOqzRsi
LHt+HtujT5c75k1lPSb9rrBtFuLYtnlzRTunsbrywl0N94XfoeZExUNqllArVnJPNx5thFgP1v2G
OvB252g8GqJB3SCTKSjVwfONGaV9J67dsoX7zuE0JGjMmoyXf9bQOmFG3MFqL22HDaMV32wREaLP
nl6YMKhvilGSbEJJ6xZxoJrNZ+NZfVqzbtyi7OYzfwX3fkZR7URer6iTAsjQoIypE7GqI82IXYlb
IP5bsLODEV+kRN6rK9Pdq/JePt4AB9NraUIj3TC8GL2nsnaSgufnK2EDz5gRtbKHfBII52gfVJ6V
GXOmuqnbNyU7+R06/3dZHuenOvK8VHbIUWVojshZEEe2ZM+i4B0AqmKWB+G2XQnnKAe9+2lU3XPF
1x7u6mstyxak7icCMwVBgQUZCLUnBAF/dQyGHrZD+yXs48f0FUBiqm5b807IiLfae1hY48K1p5cs
4N4O/G0sK03Hr++Q6XSi890iliGKuvoJyyqM8rI8jTs6gmd2VQUSxe3GixUcjOc3HL/Lui7PsngI
Cs6v4LIg5OYvLFPL7o10aa9JYFdgQ0/tO2OdGMvr2kYQNnfuIL3Yk/cDyEYWgXwS6ZBjMmYHjQI2
1pqoQv0uwYv7yulScv1ybXDa3xEGBFe4vdr9y6yTE3/KgVdkJI7lsIEunv6ryg7S6RiBjcWLDf2C
VeM9Bs5Yt6ArCnhbFtPXLjyJxZvExTjQYUdhimfoqIIZCC6cWwIHcUuoZohQGj5/dhSoeDthuPHT
kAejJ7kF+62oniTtd3WkIsl8alfngxwSOff8tY9NLqskcpwCq+juCscFSvdwZIU3lfAqS5uI6pKz
OmVcGU90sKkpPz4E21AWRYO6aTC+/lFB7RaFfVQdgf+RpVhiePrG2mNm44hO/+6tlsa8sN3N+zB5
GZMAT/5fcGhEB7tIviml7kngP2VXuNqLrxm8ZtsJiqIYyUol9KousOm6MU3AlkZPk8yZJa1pqi21
DTLUjgqCGXcY81ZkaKL3SQTPxP+DPjv8d9amMxjMOewfpy4J18JucDy/8idQHFMxyitYjQvUtx+f
xWSDrE4g9AARI9oUZI3Ez1z8jnVTKBRrAjMSaGWvxcpVUf2emSNd9h2xYkd/XArMFGvxr7GCPoLx
2VcV5sd1DG4NaUf59SSe4+hUewrLj2tV35iZtUmPN9Pq/FmYP49WWCZe+SicFa3neApA5lon09Qx
YyEZ4bkRbHIkb6Ljrgnjt9fuycuUR5tWYBzG91KN2C09hH6p2IFmg3ylku4+9X4l5lwlAWVxJd+X
KxMcRWjyitEC0TwFbzKqAtWtLETg+wvHstCSchG1iZjV/35fEBkkZVC15erlqFYDcV+bKg9uuxmi
1OIMwhodm6LkUt79ulePX+Po8qrIz5QGUlcZUJeeJf7Irsn+N9gy+x8tNalXvPSVRPbl07httINm
TqNS+gGAByWXhhTvJOc8wxzJluAPKNfsYLXsrhV7fR2Z0wpNKn3U0HnWBhGNtMmR7a+HKy+EVeGT
pH5KNLyLYI0l2UDmvqkXtgmPKDTd98j/WlLopfTDbI1pQpExP/RrRmE8qhjmtEN3yLlOjQGxdoo5
hvz2YKkra3V1tvEgv3ZhpPLkAO4L7afUHbL2EbVyGX+oFrgtXVq7GoCcdO8+88huNp8f2iXfaFyk
r/YX8Dl+MgVVscMzMrAQ3sGj9IdUQltXYMtB3eaNG3zuzuI7CZfzIczZuOwiKuXQorRl4VODXsjD
5yVWokYI2McppIglxl9bE96xVBwPfw4sbErKY/crEaFsQ1lWKYYmAO87rKMDZikcbPj/Ul5Ke4lo
DhOmjQcwByPq9GsCbAGrjcNFSQalqYgDh1ITl1k1q140c/Rbp8lxPxVgifIZsgpz7+Pq7npmA9Yt
nNUUYZvYVPwWzixzDYcLulXE3wqAKGz9MR41ao5h6vZCizluDEPs8Sp4ESmGFTPeXdZ2xDtuqLH3
dKvXeFay5L557Ysp8QYFFk/ZxA/bBUNPGnG+qOawmuHuICl2+blVOMYJcZZ9NBU4aBmSWnO+QBV/
8mrUsjE6FgMooSsTtLkS6RlMjt9S4Nxc81OiysVMFbsxolgHK03ZUi/i0NYmZWUX1j7kpWmPTdek
oJG6MCXWhg/3z6e7lDCjcSoGoz18Lrs6yWiVDWSZOUAQ07UZkt9jFLjPJzdkxgrK+5xgfe5lB3sM
gBQzZ3zrkBZPqa0dcdfQHhVV3qAO8SdHHAVXKJO5HX614Twfv3TG2Jj6YAGPLYTPPclwJExAoSwi
0GgCRYzKWsiIbQ3uT0K6297td3UBXHh0xV+Nf6rU+QrMXeLzar11R06Fj7NeTAOMloqVrgWe6V5r
nPCZlwfigexsilI9kYXDvFz36R3P/ffhIBYF0DNbiLj9FRU6LwnU5zf/nvrU0teL0vqTftYwmWgp
FlF050a0aP70LTaHzm7wAnLdyXmBHeCRKw9zH9wDmq7xdjIsP4pAUhgxQAzxq5Xb46fi80DR5u5x
A5FnHxIO+Jbxtm509SzZnpKH8h0KB5oqANvcFflforlexaJqOECR5BiCSiIfGF+65SMLYpXAmKl9
cFlRcU4X/Smaqx4TfLunMvvvbKF2uHi9wYBENmIV8dF7sTCHSbvURf+E4A9lQFzhqkhIKt+da/a0
c6gkYFL7WWDyzPetUGGkLIcf/ik921/Wlr17NmOYYfwZWmzYyBmu+TRtgbV2tU1D/Vm+Fn2NVOxd
OnbEEICtT/dRW19zQ0tL0j2pSLQ0D6y2OSug23JwAzts6so7q9/Cu13nKn2RzXxra5KNaiUFl2Oa
XIKyVZ0OjRnEzXZeX9EIAMkYuxeluX/sX28e3xxw+mVnYRrII6zWbaN63xsTJskPXqHjmT8PlW8w
86VPon/hHuqU7bDpt4tG35+zSm2Owxqwc2UV88M4f3RwFah2MFHusc6h4uXGvgzppLP7dqpHyFmK
5+OcPvGzw4ELO2E1WvfB1wWI1qFYdUYIUlbdQK9QGJsQdflVFjbzwWkKu+wvfnQPSMDCLREGsCL8
cU88++s12TLQR3Zd6u1szf0XknReAlp44YwjcANHIC/qZcXee6U4eT7Vz+QmeqbxqBm7ZJVSKGUU
mrsYCcYJBdNOx8AcPLs7PN0Qgl95N4osu0ZWOS0nVKbI/J8dqtJHYmajGriTrBwS9wn78EfWqbn7
KKIBBCox9hqU1eOflkJd4AbIemQH5jgURk8RWS6BwQpdtyn3EphiYt3zexkcLfOItMtgOu1x/nqZ
NT/9YAcUs+dA3pEPGO45uPc+KVsO+5xX66IPURDVYcf8WjDo1PyarH7hONWRgcNoXhtTxNeCoGDQ
RAy20fx+7DKIp7hj+988i8ZBDCH8/yF9TijbCwK7bX66jHgWOp5B2WzVfFk3fG8zSCTvVXaTqSjm
jtKzw8d0LiIlyvarheTe5vN/fRFTjDlYQHFHG666pbcY3AlzM1FXI4r27H7KMV+F+RWA0RQ6gT5w
8A+ReUhGDSYoAWDpnGRpLC3SdJPJwFZe1oNzLoOF3goJA8gHpQXLTxNMhiGkGft3Es4tpNndwZ+H
4o++JSc0UYMx0YRnJyH0JJPquNYH1ZueG6XzOV3l+11/AM2kvWaBSxkGco5TaErPiYKdgYc2xoPM
IGg8MEeksPS58dwkyBrfGGQhDk4q1TiOdm71qDVRmU+Pin59ZcmtGEUKnJxl5r7xnV5SBDUAwaey
DSnc+K4+HJ+3mLrlXUKrApAU9gbNTJyRja00vYutDJffMWgPHYO8CUY8xE0MRSrlKqe06HaWplIU
1TTiprx5bbdHAjA0mmK+Nr+VIctGElue+4/C64ssCDzGDs94R7BwN6iI3QwEEcsvz+MAo/GFnwkR
IHcpX/Fg+7pjjo2xRUMVcEzpmbCfs3+WSSau5I7ONygHS7HO2xEjrVWSzGTTpc1ZFXqbl1uTW94u
1tSrPB3baZtR/TMtlrfjjyci0GK1Li2wNBy13vCF+BUyFdJX6YYGTkwLqLUsM9R6mOaRV0L3jAG2
on8YemHQBBVNMBFUAEQNxO7nLlnDjEnDkFxOesdD2vQFFdDLYEn9OxmV3LoIxzPLpLWVRcz9qRw8
Nv3WuyLgb6bvgIF2151abEUT6zMh3fHBEdwp66nGkOz9xXGehT1HhgJJOsryohS6VHdwDWR2xSaB
YT5S6gBRF6R87zcLtxwvwOR5/cay9Kcvomkk59u3KbDxslPxvdlpNTP+JES3j6l1i2+4kuwsAQz3
NF0N1DGSACyXbRhDrQn8AgmgHGo0dtcSJb5C6bJYItcpnfMZ7JwloXclpU6frJbxt2kM35r3OGt1
MrGz3WvGPm24HvfIa/Of27JgWRjh98i9ItomkttZUTNU8F8oR3I7XTtjo2LfGpP9oTR0h8I/gvy/
5kkm0E7nPvCzP3wXTT3vSi7DEpk0n8e3XQnVV2BwPY/PcreiGvaVjmImP3B3JDKlIsfDeEKUum74
2bpOloiB20bDk+36qFv3SNy40ujHbdGlihKstvTsyVhPkrzdWk0/REd/FYYg7Tp9LfHxvLqS+0xX
v+ZU1mJy01kgDK332XVeaCXMdI7hsEyE8ET+eoYchqK71g6D8LCAxgIQOdqz15kzcl1WYkox2yH2
4WDWE8Pj54U2tIgO8/8hEC93X6rLbAZHduVzb50kgp7WvRR6wOPNqWU7H0UhupEEdFOzFzGDZZjE
vy+jqqx9VuaQl+iRtD1/f6f3bgdBkAY9DKKEQUGUw9I6W4YvycHsoE2wpsoHlKh6mCDCLC+HC+45
t8oPzYlp9yH9tBwtfsKrRi8p3O8QhCgKSVAUrxuUzRYtH+ERk9DOUX8sE8wGEd38WCYExkBoZXIh
d9gNaSJ6qdrqkvvuUKkCsvA8Z/ISQ8KamQVbjmTl/22//4tyzNMfp3YE34iPZxW3z8rvDvWmeCc3
rlqh6hI+PseZO1xlt4oPYO1lDTdffbWmw4MFZhLZO/z9fD4a1G9mvV2UlQ9aOb1QFBUUOkXJtDZa
mAULnlPFSvZsBmfXg5rAD9cEpIhtKYlXHklog8hs8whbQPrp3E9A0zSP3Z1aVWEuw6IqFK9DjUs3
Z1w8iUhKnrdUp1vPPP85Msjrs+FnDhaoHxGTBausA8GSM1+2yGUbEkkw130py6BFY2Mfy2VQTwC0
4FeElX5loxXXUVp1SkyU5YOsdAO8FLqWCWURqHY7wpea0RKy/avoRb3/YfVIZSwQjalU5ivCO3la
HFJQEqG3S2Du4uGWccK6108nBl1p+cGQS78dzfln3U1hN/flnoeSprvV0FnD+N9OdzREFytHGjXi
YAe6Lp1hZnuV7vK9Dw7Q0og5wGoivVR4vPINatHUMd0SLKs6vaAEhGmGsT1Uuq3PllA7c+Cmh56r
gkyZV2vdb1GEyUYVPrqmSAfBSmHu3YFMzdVogbDHsI/JAlpNL3UcpjLlDGmMgAOaY6Tk8Hbg9c/2
+vuVg9AY48BPG1hRbs9+zzLgeMyhmF+hpk7ahrZ8P23ovbGk7RDcIdmmwjVPKeFQk9fpPzQiXa5e
QCXd1V03ZPb/D0mIT/ckMtRjaWbxgJ62vM6ittu6Erq0WuqdTSiicZHZiHmY4xuDZdtz9Iv/jojj
oAi3kmBsJS2jADXzcCrVqdu2QbwU4bhKz2kFH0CxPu4sLl9IfAm1h3frChPW19xaatxZ05E8uEjj
h1y8K04bsvxQsy4GEbzqzB8jwwKEKy/oDisllt0HhS5K4wmQBtb/SHDsqVCHDmxHD6nHnX7Pryp9
HyUCnwDN7zekB2mRxYQCgJ+rLdtNMjmwAqVFORSwtSRcVMWeChmiw3K3NwnujEzRFINqIf6g6Emv
+wgiGfCr5syCuoFwAQzKARlTvD2YxF9A0TjOBRycDXC+dQFgEihoPXq7r/iW4RyLirGyhoWro8Yx
Xq9Ze5HIhFTB20F0WvvzQBMlFpjT2SMQC9tvEBKf34VJKmITxzXScQHhsDyPQl+JNJSo/iG60k/+
HDuFC5GZ1chjqcBz1oHPPxL1uvDkM28ZRvUAE3fBUaCyyTlvIEynP3d0nQVXb1mDe3AseflbSy6i
lBy80dxJYH8Ry4Hz+9YlHAPH0AlfoE0U7glNrLhNahA2BVrQDriXHTWrwGp/wThvLhGCFkpBSnDR
U06KNjvBzy3J/tFyAHjHrT9/PW8iiWc54PGwOhJRZiM4w9R9yTfhmUn5DilozBGQ/U6GmA32BmSq
BF4V1jhgzwaw4Ao5yiKf+HExGSl3KHt8d95R3iGKefKjx9+fsALD4Sska5NJ+TETPjA2MFo/Yax6
j16d2AdgZ7qCCGAr7jjwtGdBh8uQRYTEXPwDqqo4VjpnKuL1KRsEOIyjm5/Fe+QqOt3y/NUbMdN3
T48TggkjnAqkiaHmz+kXWwxqZTnbOhJc2Pp8HJEfktLeSdh98XHo5JC0IBTsjzrgbKmjeYccfqrR
UfgCiIkS70UI/5ozTVfJo/h44+2bfGFFtm2tGnXgrfLmO9yi5HgBAcp+tOhDaHdK46kZIjeCbOwC
UkxGaaBNQxdcSpV3kpnOUZlHCHqr7qsBLg2XawdAgkCaDxa4HUyplz4drDKE5ZTeSTRMwItW2wnY
RlRMc7JSwOsQTiKlTHQ6fYV/aBl92Dw3yY80JqGeNJF84ShtxAkoG6Iv8UYodHRyNhzy7dIZO+nO
7+JmTA==
`protect end_protected

